`include "/home/volplet/Escritorio/digital1v2/lab01-2024-2-garoperob/src/sum1bcc_TB.v"
`timescale 1ns/1ns
module sum1bcc (A, B, Ci,Cout,S);

  input  A;
  input  B;
  input  Ci;
  output Cout;
  output S;

  reg [1:0] st;   // REGISTRO QEU GUARDA LA SUMA 
  assign S = st[0];
  assign Cout = st[1];

  always @ ( * ) begin
  	st  = 	A+B+Ci;
  end
  
endmodule

